library verilog;
use verilog.vl_types.all;
entity ARM_datapath is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic
    );
end ARM_datapath;
