library verilog;
use verilog.vl_types.all;
entity IF_Stagr_tb is
end IF_Stagr_tb;
