library verilog;
use verilog.vl_types.all;
entity IDtb is
end IDtb;
