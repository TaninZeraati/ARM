library verilog;
use verilog.vl_types.all;
entity ConditionCheck_TB is
end ConditionCheck_TB;
