library verilog;
use verilog.vl_types.all;
entity IF_Stage_tb is
end IF_Stage_tb;
